// this module deals with all moving obstacles (i.e. cars, trains, moving railroad crossing, etc)

 
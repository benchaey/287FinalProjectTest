// This module is for all still objects / obstacles (i.e. railroad crossing posts, trees, etc) 
